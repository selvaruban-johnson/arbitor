`include "env_arbiter_transaction.sv"
`include "env_arbiter_generator.sv"
`include "env_arbiter_driver.sv"
`include "env_arbiter_interface.sv"
`include "env_arbiter_rinterface.sv"
`include "ring_counter.sv"
`include "priority_logic.sv"
`include "arbiter.sv"
`include "ring_counter_dummy.sv"
`include "priority_logic_dummy.sv"
`include "arbiter_dummy.sv"
`include "env_arbiter_coverage.sv"
`include "env_arbiter_monitor.sv"
`include "env_arbiter_scoreboard.sv"
`include "env_arbiter_environment.sv"
`include "env_arbiter_test.sv"
`include "arbiter_top.sv"