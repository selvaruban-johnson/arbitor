class env_arbiter_transaction;
rand bit ack;
rand bit [3:0] req;
bit [3:0] grant;
endclass